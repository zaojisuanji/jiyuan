----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    08:53:17 11/21/2016 
-- Design Name: 
-- Module Name:    IfIdRegisters - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity IfIdRegisters is
	--IF/ID�׶μĴ���
	port(
		rst : in std_logic;
		clk : in std_logic;
		commandIn : in std_logic_vector(15 downto 0);
		PCIn : in std_logic_vector(15 downto 0); 
		IfIdKeep : in std_logic;		--LW���ݳ�ͻ��
		IfIdFlush : in std_logic;		--��תʱ��
		
		rx : out std_logic_vector(2 downto 0);		--Command[10:8]
		ry : out std_logic_vector(2 downto 0);		--Command[7:5]
		rz : out std_logic_vector(2 downto 0);		--Command[4:2]
		imme_10_0 : out std_logic_vector(10 downto 0);	--Command[10:0]
		commandOut : out std_logic_vector(15 downto 0);
		PCOut : out std_logic_vector(15 downto 0)  --PC+1����MFPCָ���EXE��
	);
end IfIdRegisters;

architecture Behavioral of IfIdRegisters is
	signal tmpRx : std_logic_vector(2 downto 0);
	signal tmpRy : std_logic_vector(2 downto 0);
	signal tmpRz : std_logic_vector(2 downto 0);
	signal tmpImme : std_logic_vector(10 downto 0);
	signal tmpCommand : std_logic_vector(15 downto 0);
	signal tmpPC : std_logic_vector(15 downto 0);
	
begin
	rx <= tmpRx;
	ry <= tmpRy;
	rz <= tmpRz;
	imme_10_0 <= tmpImme;
	commandOut <= tmpCommand;
	PCOut <= tmpPC;
	process(rst, clk, commandIn, PCIn)
	begin 
		if (rst = '0') then	--���������źţ�ֱ������
			tmpRx 		<= (others => '0');
			tmpRy 		<= (others => '0');
			tmpRz 		<= (others => '0');
			tmpImme 		<= (others => '0');
			tmpCommand 	<= (others => '0');
			tmpPC 		<= (others => '0');
		elsif (clk'event and clk = '1') then 
			if (IfIdKeep = '0') then
				tmpRx 		<= commandIn(10 downto 8);
				tmpRy 		<= commandIn(7 downto 5);
				tmpRz 		<= commandIn(4 downto 2);
				tmpImme 		<= commandIn(10 downto 0);
				tmpCommand	<= commandIn;
				tmpPC 		<= PCIn;
			elsif (IfIdFlush <= '1') then --IfIdFlush�ò��÷���ʱ�������أ����ò��÷���IfIdKeep֮�󣿣�
				tmpRx 		<= (others => '0');
				tmpRy 		<= (others => '0');
				tmpRz 		<= (others => '0');
				tmpImme 		<= (others => '0');
				tmpCommand 	<= (others => '0');
				tmpPC 		<= (others => '0');
			end if;
		end if;
	end process;
	

end Behavioral;

